module encoder_16x4 (
    input  wire [15:0] in,
    output reg  [3:0]  out
);
    always @(*) begin
        case (in)
            16'b0000000000000001: out = 4'd0;
            16'b0000000000000010: out = 4'd1;
            16'b0000000000000100: out = 4'd2;
            16'b0000000000001000: out = 4'd3;
            16'b0000000000010000: out = 4'd4;
            16'b0000000000100000: out = 4'd5;
            16'b0000000001000000: out = 4'd6;
            16'b0000000010000000: out = 4'd7;
            16'b0000000100000000: out = 4'd8;
            16'b0000001000000000: out = 4'd9;
            16'b0000010000000000: out = 4'd10;
            16'b0000100000000000: out = 4'd11;
            16'b0001000000000000: out = 4'd12;
            16'b0010000000000000: out = 4'd13;
            16'b0100000000000000: out = 4'd14;
            16'b1000000000000000: out = 4'd15;
            default:              out = 4'bxxxx; // invalid input
        endcase
    end
endmodule